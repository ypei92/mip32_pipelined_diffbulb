library verilog;
use verilog.vl_types.all;
entity Top is
end Top;
