library verilog;
use verilog.vl_types.all;
entity ALU is
    generic(
        OP_TYPE_ALU     : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        OP_TYPE_JUMP    : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        OP_TYPE_BEQ     : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        OP_TYPE_BNE     : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        OP_TYPE_LW      : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        OP_TYPE_SW      : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        FUNC_TYPE_ADD   : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        FUNC_TYPE_SUB   : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        FUNC_TYPE_AND   : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        FUNC_TYPE_OR    : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        FUNC_TYPE_SLT   : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        FUNC_TYPE_XOR   : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        FUNC_TYPE_NOR   : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        FUNC_TYPE_ADDU  : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        FUNC_TYPE_SUBU  : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        FUNC_TYPE_SLTU  : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        FUNC_TYPE_SLL   : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        FUNC_TYPE_SRL   : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0)
    );
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        id_ex_reg_dst   : in     vl_logic;
        id_ex_alu_op    : in     vl_logic_vector(3 downto 0);
        id_ex_alu_src   : in     vl_logic;
        id_ex_mem_read  : in     vl_logic;
        id_ex_mem_write : in     vl_logic;
        id_ex_mem_to_reg: in     vl_logic;
        id_ex_reg_write : in     vl_logic;
        id_ex_branch    : in     vl_logic;
        id_ex_branch_bne: in     vl_logic;
        id_ex_reg_read_data1: in     vl_logic_vector(31 downto 0);
        id_ex_reg_read_data2: in     vl_logic_vector(31 downto 0);
        id_ex_rs        : in     vl_logic_vector(4 downto 0);
        id_ex_rt        : in     vl_logic_vector(4 downto 0);
        id_ex_rd        : in     vl_logic_vector(4 downto 0);
        id_ex_sign_extended: in     vl_logic_vector(31 downto 0);
        wb_write_data   : in     vl_logic_vector(31 downto 0);
        ex_mem_alu_result: in     vl_logic_vector(31 downto 0);
        ex_mem_rd       : in     vl_logic_vector(4 downto 0);
        mem_wb_rd       : in     vl_logic_vector(4 downto 0);
        ex_mem_reg_write_in: in     vl_logic;
        mem_wb_reg_write: in     vl_logic;
        id_ex_branch_pridictor_bit: in     vl_logic_vector(1 downto 0);
        pridictor_wrong : in     vl_logic;
        ex_mem_alu_result_out: out    vl_logic_vector(31 downto 0);
        ex_mem_reg_read_data2: out    vl_logic_vector(31 downto 0);
        ex_mem_rd_out   : out    vl_logic_vector(4 downto 0);
        ex_mem_mem_read : out    vl_logic;
        ex_mem_mem_write: out    vl_logic;
        ex_mem_mem_to_reg: out    vl_logic;
        ex_mem_reg_write: out    vl_logic;
        ex_mem_branch   : out    vl_logic;
        ex_mem_branch_bne: out    vl_logic;
        id_ex_rt_out    : out    vl_logic_vector(4 downto 0);
        id_ex_mem_read_out: out    vl_logic;
        ex_mem_branch_pridictor_bit: out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of OP_TYPE_ALU : constant is 1;
    attribute mti_svvh_generic_type of OP_TYPE_JUMP : constant is 1;
    attribute mti_svvh_generic_type of OP_TYPE_BEQ : constant is 1;
    attribute mti_svvh_generic_type of OP_TYPE_BNE : constant is 1;
    attribute mti_svvh_generic_type of OP_TYPE_LW : constant is 1;
    attribute mti_svvh_generic_type of OP_TYPE_SW : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_ADD : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_SUB : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_AND : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_OR : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_SLT : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_XOR : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_NOR : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_ADDU : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_SUBU : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_SLTU : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_SLL : constant is 1;
    attribute mti_svvh_generic_type of FUNC_TYPE_SRL : constant is 1;
end ALU;
